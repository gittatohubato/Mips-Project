
module instruction_reg ( IR, op , rs , rt , rd , first_16 ,first_26,shamt, funct );

input [31:0] IR ;
     
output reg [5:0]  op , funct ;     // 6 bits 
output reg [4:0]  rs , rt , rd , shamt ;   // 5 bits 
output reg [15:0]  first_16  ;     // 16 bits
output reg [25:0]  first_26 ;
 
always @ (IR) begin
   op <= IR[31:26];
   rs <= IR[25:21];
   rt <= IR[20:16];
   rd <= IR[15:11];
   first_16 <= IR[15:0];
   first_26 <= IR[25:0];
   funct <= IR[5:0];
   shamt <= IR[10:6];
   
end 

endmodule

