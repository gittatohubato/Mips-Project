module program_counter (clk, pcin, pcout,pcout4);

input  clk;
input [31:0] pcin;
output reg [31:0] pcout;
output reg [31:0] pcout4; 
integer flag = 0 ;     
integer file;
integer i;   

  always @(posedge clk)
      begin
if (! flag)
begin
pcout = 0 ;
flag <= 1 ;
pcout4 <= pcout + 4;
end 
       
else if(pcin<32764) 
begin 
pcout <= pcin;
pcout4 <= pcin + 4;
end

else
begin
$finish ;
$monitor ("h555h");
end

end


always @(negedge clk)
begin

if(flag)
begin
file = $fopen("C:\\Modeltech_pe_edu_10.4a\\examples\\TEXT FILE OF OUTPUTS\\PC Output Data .txt" , "a+");
$fdisplay(file,"%d\n",pcout);
$fclose(file);
end
end

endmodule


