module test(in , out);

input in;
output out;

reg[7:0] i;

i=2'b00000000;

endmodule
